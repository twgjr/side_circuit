.title KiCad schematic
V1 Net-_R1-Pad1_ 0 DC 1 
R1 Net-_R1-Pad1_ Net-_R1-Pad2_ R_US
R2 Net-_R1-Pad2_ 0 R_US
.end
